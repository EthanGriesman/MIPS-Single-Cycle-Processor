-- Ethan Griesman
-- Department of Electrical and Computer Engineering
-- Iowa State University
-- Spring 2024
--------------------------------------------------------------------------------------


-- ALU.vhd
--------------------------------------------------------------------------------------
-- DESCRIPTION: 32 bit full ALU with barrel shifter
--------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity ALU is
   port(
          inputA       : in std_logic_vector(31 downto 0); -- Operand 1
          inputB       : in std_logic_vector(31 downto 0); -- Operand 2
          i_shamt      : in std_logic_vector(4 downto 0);
          opSelect     : in std_logic_vector(3 downto 0); -- Op Select
          overflowEn   : in std_logic; 
          resultOut    : out std_logic_vector(31 downto 0); -- Result F
          overflow     : out std_logic; -- Overflow
          carryOut     : out std_logic; -- Carry out
          zeroOut      : out std_logic; -- 1 when resultOut = 0 Zero
     );
end ALU;

architecture structure of ALU is

     --AddSub
     component nbit_addsub is
     generic (N : integer := 16);
          port(i_A      : in std_logic_vector(31 downto 0);
               i_B      : in std_logic_vector(31 downto 0);
               i_AddSub : in std_logic;
               o_Sum    : out std_logic_vector(31 downto 0);
               o_Cm     : out std_logic;
               o_C      : out std_logic
          ); --Change to add previous carry as output in order to XOR for overflow
     end component;

     --barrelShift
     component barrelShifter
          port (
            iDir            : in std_logic;                       -- Right or Left shift
            iSra            : in std_logic; -- 1->signExtend 0->zeroExtend
            ishamt          : in std_logic_vector(4 downto 0);   -- Shift amount
            iInput          : in std_logic_vector(31 downto 0);  -- Input data
            oOutput         : out std_logic_vector(31 downto 0)  -- Output
          );
    end component;


    -- OR GATE --
     component org2 is
          port(i_A	: in std_logic;
               i_B	: in std_logic;
               o_F	: out std_logic);
     end component;
     
     -- AND GATE --
     component andg2 is
          port(i_A	: in std_logic;
               i_B	: in std_logic;
               o_F	: out std_logic);
     end component;
     
     -- XOR GATE -- 
     component xorg2 is
          port(i_A          : in std_logic;
               i_B          : in std_logic;
               o_F          : out std_logic);
     end component;
     
    -- One's Complement/NOT --
     component onesComp is
          generic(n: positive);
          port(
               i_D: in std_logic_vector(n-1 downto 0);
               o_O: out std_logic_vector(n-1 downto 0)
          );
     end component;


     -----------
     --Signals--
     -----------

        -- Bitwise signals --
        signal s_and                  :  std_logic_vector(31 downto 0);
        signal s_or                   :  std_logic_vector(31 downto 0);
        signal s_xor                  :  std_logic_vector(31 downto 0);
        signal s_not                  :  std_logic_vector(31 downto 0);
        signal s_nor                  :  std_logic_vector(31 downto 0);

        -- Arithmetic signals --
        signal s_sum                  :  std_logic_vector(31 downto 0);
        signal s_minus                :  std_logic;
        signal s_carry                :  std_logic;

        -- Shifter signals --
        signal s_shift                :  std_logic_vector(31 downto 0);
        signal s_sra                  :  std_logic_vector(31 downto 0);
        signal s_dir                  :  std_logic_vector(31 downto 0);
        signal s_shamt                :  std_logic_vector(31 downto 0);

        -- Misc signals --    
        signal s_slt                  :  std_logic_vector(31 downto 0);
        signal s_sltSum               :  std_logic_vector(31 downto 0);
        signal s_sltC                 :  std_logic_vector(31 downto 0);
        signal s_sltOverflow          :  std_logic_vector(31 downto 0);
        signal s_sltOverflowCheck     :  std_logic_vector(31 downto 0);

        -- ALU signal
        signal s_resultout            :  std_logic_vector(31 downto 0);
        signal s_zero                 :  std_logic;

        -- Overflow signal --
        signal s_overflowCheck        :  std_logic_vector(3 downto 0);
        signal s_overflow             :  std_logic;



        signal s_sll                  :  std_logic_vector(31 downto 0);
        signal s_srl                  :  std_logic_vector(31 downto 0);
        signal s_sra                  :  std_logic_vector(31 downto 0);
        signal s_sllv                 :  std_logic_vector(31 downto 0);
        signal s_srlv                 :  std_logic_vector(31 downto 0);
        signal s_srav                 :  std_logic_vector(31 downto 0);
        signal s_lui                  :  std_logic_vector(31 downto 0);

        
        begin

          -- AND --
          ALU_AND: for i in 0 to 31 generate
           ANDGS: andg2
           port map(i_A => inputA(i),
                    i_B => inputB(i),
                    o_F => s_and(i));
          end generate ALU_AND;

          -- OR --
          ALU_OR: for i in 0 to 31 generate
           ORGS: org2
           port map(i_A => inputA(i),
                    i_B => inputB(i), 
                    o_F => s_or(i));
          end generate ALU_OR;


          -- XOR --
          ALU_XOR: for i in 0 to 31 generate
           XORGS: xorg2
           port map(i_A => inputA(i),
                    i_B => inputB(i),
                    o_F => s_xor(i));
          end generate ALU_XOR;
          
          -- NOR --
          ALU_NOR: onesComp
          generic map (32)
          port map(i_D => s_or,
                   o_O => s_nor);

          -- NOT --
          ALU_NOT: onesComp
          generic map(32)
          port map(i_D => inputA,
                   o_O => s_not);

          
          -- ADD SUB --
          adderN : n_addsub
           port map(iA => inputA,
                    iB => inputB,
                    i_AddSub => s_minus,       -- 
                    iC => i_Op(0),   -- carry in 
                    oC => s_carry,    -- carry out
                    oS => s_sum); -- sum output


          -- 0 for left, 1 for right --          
          with opSelect select 
            s_dir <= '0' when "1000" | "1011"
                     '1' when others;
          
          -- 0 for logical, 1 for arithmetic --
          with opSelect select 
            s_sra <= '0' when "1000" | "1011"
                     '1' when others;
         
          with opSelect select 
            s_shamt <= i_shamt when "1000" | "1001" | "1010",
                      when others;

          -- Barrel Shifter
          ALU_SHIFTER: barrelShifter
           generic map(32)
           port map(
                    iInput  => inputB,
                    i_shamt => s_shamt,
                    iDir => s_dir,  -- Perform subtraction: inputA - inputB
                    iSra => s_sra,  -- The subtraction result
                    o_C => s_shift       -- Ignore carry-out
               );

          -- SLT
          s_sltOverflowCheck <= i_Ain(31) & i_Bin(31) & s_sltSum(31);
          with s_sltOverflowCheck select
            s_sltOverflowCheck <= '1' when "001",
                                  '1' when "100",
                                  '1' when "101",
                                  '1' when "111",
                                  '0' when others;

          ALU_SLT: n_addsub
          port map(i_A => inputA,
                    i_B => inputB,
                    i_AddSub => '1',       -- 
                    iC => i_Op(0),   -- carry in 
                    oC => s_sltSum,    -- carry out
                    oS => s_sltC); -- sum output


          -- signal is 1 or 0
          s_slt <= "0000000000000000000000000000000" & s_sltOverflow;
          
          -- LUI --
          s_lui <= inputB(15 downto 0)&"0000000000000000";


          --Output Selection--
          with opSelect select  --diff than add sub
          s_resultout <= s_add when "000000000", --add/sub  
                         s_and when "000000011", --and
                         s_nor when "000010010", --nor
                         s_xor when "000000100", --xor
                         s_or when "000000010", --or
                         s_slt when "100000101", --slt
                         --s_sll when "000000001" , --sll
                         --s_srl when "000001001", --srl
                         --s_sra when "010001001", --sra
                         s_sub when "100000000", --sub
                         -- s_sllv when "000100001", --sllv
                         -- s_srlv when "000101001", --srlv
                         -- s_srav when "010101001", --srav
                         -- s_lui when "001000001", --lui
                         "11111111111111111111111111111111" when others;

          with s_resultout select
            s_zero <= '1' when "0000000000000000000000000000000",
                      '0' when others;

          o_aluOut <= s_aluOut;
          o_zero <= s_zero;
          o_carry <= s_carry;

          -- Logic for overflow
          s_overflowCheck <= inputA(31) & inputB(31) & s_minus & s_sum(31);
          with s_overflowCHeck select
            s_overflow <= '1' when "001",
                                  '1' when "0001",
                                  '1' when "1100",
                                  '1' when "0111",
                                  '1' when "1010",
                                  '0' when others;

          overflow <= s_overflow AND overflowEn;

end structure;
        
    